`timescale 1ns / 100ps
// nano = 10^-9
// pico = 10^-12
// Timescale specifies the time unit and time precision 
// of a module that follow it. The simulation time and delay
// values are measured using time unit. The precision factor
// is needed to measure the degree of accuracy of the time
// unit, in other words how delay values are rounded before
// being used in simulation.
